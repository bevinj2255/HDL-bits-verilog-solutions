module top_module(input in, output wire out );
    assign out = in;
endmodule
